/* Control Unit */

`timescale 1ns/1ns

`ifndef _datapath
`define _datapath

module datapath(
  
);


endmodule

`endif