/* 4 to 16 demultiplexer (decoder) */

`timescale 1ns/1ns

module dmux4x16(
  input  en,
  input  [3:0] sel,
  output reg [15:0] d
);

  always @(sel or en) begin
    d = 16'b0;
    if(en) begin
      case(sel)
        4'b0000: d = 16'b0000000000000001; // R0
        4'b0001: d = 16'b0000000000000010; // R1
        4'b0010: d = 16'b0000000000000100; // R2
        4'b0011: d = 16'b0000000000001000; // R3
        4'b0100: d = 16'b0000000000010000; // R4
        4'b0101: d = 16'b0000000000100000; // R5
        4'b0110: d = 16'b0000000001000000; // R6
        4'b0111: d = 16'b0000000010000000; // R7
        4'b1000: d = 16'b0000000100000000; // R8
        4'b1001: d = 16'b0000001000000000; // R9
        4'b1010: d = 16'b0000010000000000; // R10
        4'b1011: d = 16'b0000100000000000; // R11
        4'b1100: d = 16'b0001000000000000; // R12
        4'b1101: d = 16'b0010000000000000; // R13
        4'b1110: d = 16'b0100000000000000; // R14
        4'b1111: d = 16'b1000000000000000; // R15
        default: d = 16'b0000000000000000; // invalid state
      endcase
    end
  end

endmodule