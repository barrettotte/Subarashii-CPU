/* Control Unit */

`timescale 1ns/1ns

`ifndef _cu
`define _cu

module cu(
  
);



endmodule

`endif